library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 8;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
        -- Inicializa os endereços:
tmp(0) := x"9" & "00" & '0' & x"24";	-- JSR .setup          	# Chama a função setup, para limpar os endereços
tmp(1) := x"6" & "00" & '0' & x"07";	-- JMP .LOOP_HEX
tmp(2) := x"9" & "00" & '0' & x"B3";	-- JSR .troca_hex PASSA_HEX:          # começo do LOOP para HEX0
tmp(3) := x"6" & "00" & '0' & x"07";	-- JMP .LOOP_HEX
tmp(4) := x"9" & "00" & '0' & x"B0";	-- JSR .limpa_but VOLTA_SET_RELOGIO:
tmp(5) := x"9" & "00" & '1' & x"7C";	-- JSR .setar_hora
tmp(6) := x"9" & "00" & '1' & x"55";	-- JSR .ajusta_leds
tmp(7) := x"9" & "00" & '0' & x"4A";	-- JSR .logica_seleciona LOOP_HEX:
tmp(8) := x"7" & "00" & '0' & x"02";	-- JEQ .PASSA_HEX       	# SE botão for pressionado realiza o salto, se não continua
tmp(9) := x"9" & "00" & '0' & x"52";	-- JSR .verifica_key1
tmp(10) := x"7" & "00" & '0' & x"0C";	-- JEQ .relogio_principal
tmp(11) := x"6" & "00" & '0' & x"07";	-- JMP .LOOP_HEX      	# se botão não pressionado, volta para o LOOP de HEX0
tmp(12) := x"9" & "00" & '0' & x"B0";	-- JSR .limpa_but relogio_principal:
tmp(13) := x"9" & "00" & '1' & x"79";	-- JSR .limpa_led
tmp(14) := x"9" & "00" & '0' & x"4E";	-- JSR .verifica_key0 loop_relogio:
tmp(15) := x"7" & "00" & '0' & x"04";	-- JEQ .VOLTA_SET_RELOGIO
tmp(16) := x"9" & "00" & '0' & x"C3";	-- JSR .verifica_carry
tmp(17) := x"1" & "10" & '1' & x"62";	-- LDA R2 @KEY2
tmp(18) := x"8" & "10" & '0' & x"00";	-- CEQ R2 @ZERO
tmp(19) := x"7" & "00" & '0' & x"19";	-- JEQ .TEMPO_RAPIDO
tmp(20) := x"4" & "11" & '0' & x"00";	-- LDI R3 $0
tmp(21) := x"5" & "11" & '1' & x"00";	-- STA @LED0A7 R3
tmp(22) := x"1" & "00" & '1' & x"65";	-- LDA R0 @BASE_TEMPO        		# Salva o endereço da base_tempo2 no R0
tmp(23) := x"5" & "00" & '1' & x"FD";	-- STA @LIMPA_BASE_TEMPO R0    
tmp(24) := x"6" & "00" & '0' & x"1D";	-- JMP .VERIFICA_TEMPO
tmp(25) := x"4" & "11" & '0' & x"40";	-- LDI R3 $64 TEMPO_RAPIDO:
tmp(26) := x"5" & "11" & '1' & x"00";	-- STA @LED0A7 R3
tmp(27) := x"1" & "00" & '1' & x"66";	-- LDA R0 @BASE_TEMPO_RAP        		# Salva o endereço da base_tempo2 no R0
tmp(28) := x"5" & "00" & '1' & x"FC";	-- STA @LIMPA_BASE_TEMPO_RAP R0  
tmp(29) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM                  	# Verifica se a base de tempo será utilizada VERIFICA_TEMPO:
tmp(30) := x"7" & "00" & '0' & x"20";	-- JEQ .INCREMENTA             	# Se for vai para a rotina de incremento
tmp(31) := x"6" & "00" & '0' & x"0E";	-- JMP .loop_relogio
tmp(32) := x"1" & "01" & '0' & x"14";	-- LDA R1 @VALOR_ATUAL0 INCREMENTA:
tmp(33) := x"2" & "01" & '0' & x"01";	-- SOMA R1 @UM
tmp(34) := x"5" & "01" & '0' & x"14";	-- STA @VALOR_ATUAL0 R1
tmp(35) := x"6" & "00" & '0' & x"0E";	-- JMP .loop_relogio
tmp(36) := x"0" & "00" & '0' & x"00";	-- NOP setup:              # Definindo a função setup, roda sempre no início limpando os valores
tmp(37) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0           
tmp(38) := x"5" & "00" & '0' & x"00";	-- STA @ZERO R0
tmp(39) := x"5" & "00" & '0' & x"06";	-- STA @ATUAL R0
tmp(40) := x"5" & "00" & '1' & x"20";	-- STA @HEX0 R0
tmp(41) := x"5" & "00" & '1' & x"21";	-- STA @HEX1 R0
tmp(42) := x"5" & "00" & '1' & x"22";	-- STA @HEX2 R0
tmp(43) := x"5" & "00" & '1' & x"23";	-- STA @HEX3 R0
tmp(44) := x"5" & "00" & '1' & x"24";	-- STA @HEX4 R0
tmp(45) := x"5" & "00" & '1' & x"25";	-- STA @HEX5 R0
tmp(46) := x"5" & "00" & '1' & x"01";	-- STA @LED8 R0
tmp(47) := x"5" & "00" & '1' & x"02";	-- STA @LED9 R0
tmp(48) := x"5" & "00" & '0' & x"14";	-- STA @VALOR_ATUAL0 R0
tmp(49) := x"5" & "00" & '0' & x"15";	-- STA @VALOR_ATUAL1 R0
tmp(50) := x"5" & "00" & '0' & x"16";	-- STA @VALOR_ATUAL2 R0
tmp(51) := x"5" & "00" & '0' & x"17";	-- STA @VALOR_ATUAL3 R0
tmp(52) := x"5" & "00" & '0' & x"18";	-- STA @VALOR_ATUAL4 R0
tmp(53) := x"5" & "00" & '0' & x"19";	-- STA @VALOR_ATUAL5 R0
tmp(54) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1
tmp(55) := x"5" & "00" & '0' & x"01";	-- STA @UM R0
tmp(56) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(57) := x"5" & "00" & '1' & x"FF";	-- STA @LIMPA_KEY0 R0
tmp(58) := x"4" & "00" & '0' & x"02";	-- LDI R0 $2
tmp(59) := x"5" & "00" & '0' & x"02";	-- STA @DOIS R0
tmp(60) := x"4" & "00" & '0' & x"03";	-- LDI R0 $3
tmp(61) := x"5" & "00" & '0' & x"03";	-- STA @TRES R0
tmp(62) := x"4" & "00" & '0' & x"04";	-- LDI R0 $4
tmp(63) := x"5" & "00" & '0' & x"04";	-- STA @QUATRO R0
tmp(64) := x"4" & "00" & '0' & x"05";	-- LDI R0 $5
tmp(65) := x"5" & "00" & '0' & x"05";	-- STA @CINCO R0
tmp(66) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(67) := x"4" & "00" & '0' & x"06";	-- LDI R0 $6
tmp(68) := x"5" & "00" & '0' & x"25";	-- STA @SEIS R0
tmp(69) := x"4" & "00" & '0' & x"0A";	-- LDI R0 $10
tmp(70) := x"5" & "00" & '0' & x"26";	-- STA @DEZ R0
tmp(71) := x"4" & "00" & '0' & x"20";	-- LDI R0 $32
tmp(72) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(73) := x"A" & "00" & '0' & x"00";	-- RET
tmp(74) := x"9" & "00" & '0' & x"56";	-- JSR .escreveSW      	# Função que realiza a leitura e faz verificação em qual HEX está escrevendo e escreve no correto logica_seleciona:
tmp(75) := x"9" & "00" & '0' & x"B7";	-- JSR .verifica_SW9   	# Função que faz a verificação se o SW9 está ativo, se sim será 12H
tmp(76) := x"9" & "00" & '0' & x"4E";	-- JSR .verifica_key0  	# Função que faz a verificação se o botão KEY0 foi pressionado, se sim flag EQUAL = 1
tmp(77) := x"A" & "00" & '0' & x"00";	-- RET
tmp(78) := x"0" & "00" & '0' & x"00";	-- NOP verifica_key0:      # Definindo a função para verificar KEY0
tmp(79) := x"1" & "10" & '1' & x"60";	-- LDA R2 @KEY0
tmp(80) := x"8" & "10" & '0' & x"01";	-- CEQ R2 @UM
tmp(81) := x"A" & "00" & '0' & x"00";	-- RET
tmp(82) := x"0" & "00" & '0' & x"00";	-- NOP verifica_key1:      # Definindo a função para verificar KEY1
tmp(83) := x"1" & "11" & '1' & x"61";	-- LDA R3 @KEY1
tmp(84) := x"8" & "11" & '0' & x"01";	-- CEQ R3 @UM
tmp(85) := x"A" & "00" & '0' & x"00";	-- RET
tmp(86) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7 escreveSW:
tmp(87) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(88) := x"8" & "00" & '0' & x"05";	-- CEQ R0 @CINCO
tmp(89) := x"7" & "00" & '0' & x"9A";	-- JEQ .HEX5 
tmp(90) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(91) := x"8" & "00" & '0' & x"04";	-- CEQ R0 @QUATRO
tmp(92) := x"7" & "00" & '0' & x"81";	-- JEQ .HEX4
tmp(93) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(94) := x"8" & "00" & '0' & x"03";	-- CEQ R0 @TRES
tmp(95) := x"7" & "00" & '0' & x"7B";	-- JEQ .HEX3 
tmp(96) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(97) := x"8" & "00" & '0' & x"02";	-- CEQ R0 @DOIS
tmp(98) := x"7" & "00" & '0' & x"75";	-- JEQ .HEX2
tmp(99) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(100) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(101) := x"7" & "00" & '0' & x"6F";	-- JEQ .HEX1
tmp(102) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(103) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(104) := x"7" & "00" & '0' & x"69";	-- JEQ .HEX0
tmp(105) := x"C" & "01" & '0' & x"26";	-- CLT R1 @DEZ HEX0:
tmp(106) := x"D" & "00" & '0' & x"6C";	-- JLT .CARREGA_HEX0
tmp(107) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(108) := x"5" & "01" & '1' & x"20";	-- STA @HEX0 R1 CARREGA_HEX0:
tmp(109) := x"5" & "01" & '0' & x"14";	-- STA @VALOR_ATUAL0 R1 
tmp(110) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL 
tmp(111) := x"C" & "01" & '0' & x"25";	-- CLT R1 @SEIS  HEX1:
tmp(112) := x"D" & "00" & '0' & x"72";	-- JLT .CARREGA_HEX1
tmp(113) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(114) := x"5" & "01" & '1' & x"21";	-- STA @HEX1 R1  CARREGA_HEX1:
tmp(115) := x"5" & "01" & '0' & x"15";	-- STA @VALOR_ATUAL1 R1 
tmp(116) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL 
tmp(117) := x"C" & "01" & '0' & x"26";	-- CLT R1 @DEZ HEX2:
tmp(118) := x"D" & "00" & '0' & x"78";	-- JLT .CARREGA_HEX2
tmp(119) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(120) := x"5" & "01" & '1' & x"22";	-- STA @HEX2 R1  CARREGA_HEX2:
tmp(121) := x"5" & "01" & '0' & x"16";	-- STA @VALOR_ATUAL2 R1 
tmp(122) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL 
tmp(123) := x"C" & "01" & '0' & x"25";	-- CLT R1 @SEIS HEX3:
tmp(124) := x"D" & "00" & '0' & x"7E";	-- JLT .CARREGA_HEX3
tmp(125) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(126) := x"5" & "01" & '1' & x"23";	-- STA @HEX3 R1  CARREGA_HEX3:
tmp(127) := x"5" & "01" & '0' & x"17";	-- STA @VALOR_ATUAL3 R1 
tmp(128) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL 
tmp(129) := x"1" & "00" & '0' & x"1F";	-- LDA R0 @FLAG_12_OU_24 HEX4:
tmp(130) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(131) := x"7" & "00" & '0' & x"8E";	-- JEQ .12_VERIFICA
tmp(132) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5
tmp(133) := x"8" & "10" & '0' & x"02";	-- CEQ R2 @DOIS 
tmp(134) := x"7" & "00" & '0' & x"8A";	-- JEQ .HEX5_DOIS
tmp(135) := x"C" & "01" & '0' & x"26";	-- CLT R1 @DEZ 
tmp(136) := x"D" & "00" & '0' & x"97";	-- JLT .CARREGA_HEX4
tmp(137) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(138) := x"C" & "01" & '0' & x"04";	-- CLT R1 @QUATRO  HEX5_DOIS:
tmp(139) := x"D" & "00" & '0' & x"97";	-- JLT .CARREGA_HEX4 
tmp(140) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(141) := x"7" & "00" & '0' & x"97";	-- JEQ .CARREGA_HEX4
tmp(142) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5 12_VERIFICA:
tmp(143) := x"8" & "10" & '0' & x"00";	-- CEQ R2 @ZERO 
tmp(144) := x"7" & "00" & '0' & x"94";	-- JEQ .12_HEX5_ZERO
tmp(145) := x"C" & "01" & '0' & x"03";	-- CLT R1 @TRES
tmp(146) := x"D" & "00" & '0' & x"97";	-- JLT .CARREGA_HEX4
tmp(147) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(148) := x"C" & "01" & '0' & x"26";	-- CLT R1 @DEZ 12_HEX5_ZERO:
tmp(149) := x"D" & "00" & '0' & x"97";	-- JLT .CARREGA_HEX4
tmp(150) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(151) := x"5" & "01" & '1' & x"24";	-- STA @HEX4 R1  CARREGA_HEX4:
tmp(152) := x"5" & "01" & '0' & x"18";	-- STA @VALOR_ATUAL4 R1 
tmp(153) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL 
tmp(154) := x"1" & "00" & '0' & x"1F";	-- LDA R0 @FLAG_12_OU_24           	# Verifica se está no modo 12H ou 24H HEX5:
tmp(155) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM                      	# Se estiver no modo de 12H ele salta
tmp(156) := x"7" & "00" & '0' & x"A0";	-- JEQ .12_VERIFICA_5              	# Salta se 12H estiver ativado
tmp(157) := x"C" & "01" & '0' & x"03";	-- CLT R1 @TRES                    	# Se estiver no modo 24H verifica a flag para ver se é menor que 3
tmp(158) := x"D" & "00" & '0' & x"A3";	-- JLT .CARREGA_HEX5
tmp(159) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(160) := x"C" & "01" & '0' & x"02";	-- CLT R1 @DOIS                   	# Verifica a flag_1, que ativa se o valor dos SW for menor que 2 12_VERIFICA_5:
tmp(161) := x"D" & "00" & '0' & x"A3";	-- JLT .CARREGA_HEX5
tmp(162) := x"6" & "00" & '0' & x"A5";	-- JMP .FINAL
tmp(163) := x"5" & "01" & '1' & x"25";	-- STA @HEX5 R1  CARREGA_HEX5:                   # Escreve no HEX5
tmp(164) := x"5" & "01" & '0' & x"19";	-- STA @VALOR_ATUAL5 R1 
tmp(165) := x"A" & "00" & '0' & x"00";	-- RET  FINAL:
tmp(166) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED atualiza_atual:
tmp(167) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(168) := x"7" & "00" & '0' & x"AD";	-- JEQ .VOLTA_CINCO
tmp(169) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(170) := x"3" & "00" & '0' & x"01";	-- SUB R0 @UM
tmp(171) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(172) := x"A" & "00" & '0' & x"00";	-- RET
tmp(173) := x"4" & "00" & '0' & x"05";	-- LDI R0 $5 VOLTA_CINCO:
tmp(174) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(175) := x"A" & "00" & '0' & x"00";	-- RET
tmp(176) := x"5" & "00" & '1' & x"FF";	-- STA @LIMPA_KEY0 R0  limpa_but:
tmp(177) := x"5" & "00" & '1' & x"FE";	-- STA @LIMPA_KEY1 R0
tmp(178) := x"A" & "00" & '0' & x"00";	-- RET
tmp(179) := x"9" & "00" & '0' & x"A6";	-- JSR .atualiza_atual troca_hex:
tmp(180) := x"9" & "00" & '1' & x"55";	-- JSR .ajusta_leds
tmp(181) := x"9" & "00" & '0' & x"B0";	-- JSR .limpa_but
tmp(182) := x"A" & "00" & '0' & x"00";	-- RET
tmp(183) := x"1" & "00" & '1' & x"42";	-- LDA R0 @SW9 verifica_SW9:
tmp(184) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(185) := x"7" & "00" & '0' & x"BE";	-- JEQ .SW_ATIVO
tmp(186) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(187) := x"5" & "00" & '0' & x"1F";	-- STA @FLAG_12_OU_24 R0 
tmp(188) := x"5" & "00" & '1' & x"02";	-- STA @LED9 R0
tmp(189) := x"A" & "00" & '0' & x"00";	-- RET
tmp(190) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1 SW_ATIVO:
tmp(191) := x"5" & "00" & '0' & x"1F";	-- STA @FLAG_12_OU_24 R0 
tmp(192) := x"5" & "00" & '1' & x"02";	-- STA @LED9 R0
tmp(193) := x"9" & "00" & '1' & x"7F";	-- JSR .AM_PM
tmp(194) := x"A" & "00" & '0' & x"00";	-- RET
tmp(195) := x"1" & "10" & '0' & x"14";	-- LDA R2 @VALOR_ATUAL0            	# LEITURA DE HEX0  verifica_carry:
tmp(196) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ                     	# VERIFICA SE É IGUAL A 10 PARA O CARRY
tmp(197) := x"7" & "00" & '0' & x"C9";	-- JEQ .CARRY_DEZ_SEG              	# SALTA SE TIVER O CARRY
tmp(198) := x"1" & "10" & '0' & x"14";	-- LDA R2 @VALOR_ATUAL0            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX0
tmp(199) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(200) := x"A" & "00" & '0' & x"00";	-- RET
tmp(201) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO                    	# COMO TEVE O CARRY, ESCREVE 0 EM SEGUNDO CARRY_DEZ_SEG:
tmp(202) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(203) := x"5" & "10" & '0' & x"14";	-- STA @VALOR_ATUAL0 R2        	# ESCREVE 0 NOS SEGUNDOS QUANDO CARRY
tmp(204) := x"1" & "10" & '0' & x"15";	-- LDA R2 @VALOR_ATUAL1        	# LEITURA DO HEX1
tmp(205) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(206) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2
tmp(207) := x"8" & "10" & '0' & x"25";	-- CEQ R2 @SEIS                	# VERIFICA SE NÃO VAI TER O CARRY
tmp(208) := x"7" & "00" & '0' & x"D4";	-- JEQ .CARRY_MIN              	# SALTA SE TIVER CARRY
tmp(209) := x"1" & "10" & '0' & x"15";	-- LDA R2 @VALOR_ATUAL1            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX1
tmp(210) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(211) := x"A" & "00" & '0' & x"00";	-- RET
tmp(212) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO                	# COMO TEVE CARRY ESCREVE 0 EM HEX1 CARRY_MIN:
tmp(213) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(214) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2 
tmp(215) := x"1" & "10" & '0' & x"16";	-- LDA R2 @VALOR_ATUAL2        	# LEITURA DO HEX2 PARA VER SE VAI TER CARRY
tmp(216) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(217) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2
tmp(218) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ
tmp(219) := x"7" & "00" & '0' & x"DF";	-- JEQ .CARRY_DEZ_MIN          	# SE TIVER CARRY REALIZA O SALTO
tmp(220) := x"1" & "10" & '0' & x"16";	-- LDA R2 @VALOR_ATUAL2            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX2
tmp(221) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(222) := x"A" & "00" & '0' & x"00";	-- RET
tmp(223) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO               	# COMO TEVE CARRY ESCREVE 0 EM HEX2 CARRY_DEZ_MIN:
tmp(224) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(225) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2 
tmp(226) := x"1" & "10" & '0' & x"17";	-- LDA R2 @VALOR_ATUAL3
tmp(227) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(228) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2
tmp(229) := x"8" & "10" & '0' & x"25";	-- CEQ R2 @SEIS
tmp(230) := x"7" & "00" & '0' & x"EA";	-- JEQ .CARRY_HORA
tmp(231) := x"1" & "10" & '0' & x"17";	-- LDA R2 @VALOR_ATUAL3            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX3
tmp(232) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(233) := x"A" & "00" & '0' & x"00";	-- RET
tmp(234) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO CARRY_HORA:
tmp(235) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(236) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2 
tmp(237) := x"1" & "11" & '0' & x"1F";	-- LDA R3 @FLAG_12_OU_24
tmp(238) := x"8" & "11" & '0' & x"01";	-- CEQ R3 @UM
tmp(239) := x"7" & "00" & '1' & x"1E";	-- JEQ .HORA_12        	#SALTA SE O MODO DE 12 HORAS ESTIVER ATIVADO 
tmp(240) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4        	# COMEÇA A VERIFICAÇÃO PARA 24HORAS
tmp(241) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(242) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(243) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5        	# PEGA O VALOR DA HORA PARA SABER QUAL COMPARAÇÃO VOCÊ VAI FAZER
tmp(244) := x"8" & "10" & '0' & x"02";	-- CEQ R2 @DOIS 
tmp(245) := x"7" & "00" & '0' & x"FC";	-- JEQ .DEPOIS_DAS_20H
tmp(246) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(247) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ
tmp(248) := x"7" & "00" & '1' & x"16";	-- JEQ .CARRY_HORA_24
tmp(249) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX2
tmp(250) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(251) := x"A" & "00" & '0' & x"00";	-- RET                           	# ROTINA ANTES DAS 20H
tmp(252) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4 DEPOIS_DAS_20H:
tmp(253) := x"8" & "10" & '0' & x"04";	-- CEQ R2 @QUATRO 
tmp(254) := x"7" & "00" & '1' & x"08";	-- JEQ .RESET_24_HORA
tmp(255) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(256) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2 
tmp(257) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(258) := x"A" & "00" & '0' & x"00";	-- RET
tmp(259) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	#QUANDO ESTAMOS EM 20HORAS MAIS
tmp(260) := x"8" & "10" & '0' & x"04";	-- CEQ R2 @QUATRO
tmp(261) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX4 JEQ .RESET_24_HORA:
tmp(262) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(263) := x"A" & "00" & '0' & x"00";	-- RET
tmp(264) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO RESET_24_HORA:
tmp(265) := x"5" & "10" & '0' & x"14";	-- STA @VALOR_ATUAL0 R2 
tmp(266) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(267) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2 
tmp(268) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(269) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2 
tmp(270) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(271) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2
tmp(272) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(273) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(274) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(275) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(276) := x"5" & "10" & '1' & x"25";	-- STA @HEX5 R2
tmp(277) := x"A" & "00" & '0' & x"00";	-- RET
tmp(278) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO CARRY_HORA_24:
tmp(279) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(280) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2 
tmp(281) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5
tmp(282) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(283) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(284) := x"5" & "10" & '1' & x"25";	-- STA @ HEX5 R2
tmp(285) := x"A" & "00" & '0' & x"00";	-- RET
tmp(286) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4        	# LEITURA DE HEX4 HORA_12:
tmp(287) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(288) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(289) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5
tmp(290) := x"8" & "10" & '0' & x"01";	-- CEQ R2 @UM
tmp(291) := x"7" & "00" & '1' & x"2A";	-- JEQ .10H_MAIS
tmp(292) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(293) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ
tmp(294) := x"7" & "00" & '1' & x"34";	-- JEQ .CARRY_DEZ_HORA_12
tmp(295) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(296) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(297) := x"A" & "00" & '0' & x"00";	-- RET 
tmp(298) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4 10H_MAIS:
tmp(299) := x"8" & "10" & '0' & x"03";	-- CEQ R2 @TRES
tmp(300) := x"7" & "00" & '1' & x"3C";	-- JEQ .RESET_12H_TROCA_AM_PM
tmp(301) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(302) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(303) := x"A" & "00" & '0' & x"00";	-- RET 
tmp(304) := x"7" & "00" & '1' & x"34";	-- JEQ .CARRY_DEZ_HORA_12
tmp(305) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX2
tmp(306) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(307) := x"A" & "00" & '0' & x"00";	-- RET
tmp(308) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO CARRY_DEZ_HORA_12:
tmp(309) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2 
tmp(310) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(311) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5
tmp(312) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(313) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(314) := x"5" & "10" & '1' & x"25";	-- STA @HEX5 R2
tmp(315) := x"A" & "00" & '0' & x"00";	-- RET
tmp(316) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO RESET_12H_TROCA_AM_PM:
tmp(317) := x"5" & "10" & '0' & x"14";	-- STA @VALOR_ATUAL0 R2 
tmp(318) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(319) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2 
tmp(320) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(321) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2 
tmp(322) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(323) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2
tmp(324) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(325) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(326) := x"5" & "10" & '1' & x"25";	-- STA @HEX5 R2
tmp(327) := x"1" & "10" & '0' & x"01";	-- LDA R2 @UM 
tmp(328) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(329) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(330) := x"1" & "10" & '0' & x"07";	-- LDA R2 @TROCA_AM_PM
tmp(331) := x"8" & "10" & '0' & x"00";	-- CEQ R2 @ZERO
tmp(332) := x"7" & "00" & '1' & x"51";	-- JEQ .LED8_ZERO
tmp(333) := x"1" & "10" & '0' & x"00";	-- LDA R2 $0
tmp(334) := x"5" & "10" & '1' & x"01";	-- STA @LED8 R2
tmp(335) := x"5" & "10" & '0' & x"07";	-- STA @TROCA_AM_PM R2
tmp(336) := x"6" & "00" & '1' & x"54";	-- JMP .FIM_RESET_LED8
tmp(337) := x"4" & "10" & '0' & x"01";	-- LDI R2 $1 LED8_ZERO:
tmp(338) := x"5" & "10" & '1' & x"01";	-- STA @LED8 R2
tmp(339) := x"5" & "10" & '0' & x"07";	-- STA @TROCA_AM_PM R2
tmp(340) := x"A" & "00" & '0' & x"00";	-- RET FIM_RESET_LED8:
tmp(341) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED ajusta_leds:
tmp(342) := x"8" & "00" & '0' & x"05";	-- CEQ R0 @CINCO
tmp(343) := x"7" & "00" & '1' & x"67";	-- JEQ .32_NO_LED
tmp(344) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(345) := x"8" & "00" & '0' & x"04";	-- CEQ R0 @QUATRO
tmp(346) := x"7" & "00" & '1' & x"6A";	-- JEQ .16_NO_LED
tmp(347) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(348) := x"8" & "00" & '0' & x"03";	-- CEQ R0 @TRES
tmp(349) := x"7" & "00" & '1' & x"6D";	-- JEQ .8_NO_LED
tmp(350) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(351) := x"8" & "00" & '0' & x"02";	-- CEQ R0 @DOIS
tmp(352) := x"7" & "00" & '1' & x"70";	-- JEQ .4_NO_LED
tmp(353) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(354) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(355) := x"7" & "00" & '1' & x"73";	-- JEQ .2_NO_LED
tmp(356) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(357) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(358) := x"7" & "00" & '1' & x"76";	-- JEQ .1_NO_LED
tmp(359) := x"4" & "00" & '0' & x"20";	-- LDI R0 $32 32_NO_LED:
tmp(360) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(361) := x"A" & "00" & '0' & x"00";	-- RET
tmp(362) := x"4" & "00" & '0' & x"10";	-- LDI R0 $16 16_NO_LED:
tmp(363) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(364) := x"A" & "00" & '0' & x"00";	-- RET
tmp(365) := x"4" & "00" & '0' & x"08";	-- LDI R0 $8 8_NO_LED:
tmp(366) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(367) := x"A" & "00" & '0' & x"00";	-- RET
tmp(368) := x"4" & "00" & '0' & x"04";	-- LDI R0 $4 4_NO_LED:
tmp(369) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(370) := x"A" & "00" & '0' & x"00";	-- RET
tmp(371) := x"4" & "00" & '0' & x"02";	-- LDI R0 $2 2_NO_LED:
tmp(372) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(373) := x"A" & "00" & '0' & x"00";	-- RET
tmp(374) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1 1_NO_LED:
tmp(375) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(376) := x"A" & "00" & '0' & x"00";	-- RET 
tmp(377) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0 limpa_led:
tmp(378) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(379) := x"A" & "00" & '0' & x"00";	-- RET
tmp(380) := x"4" & "00" & '0' & x"05";	-- LDI R0 $5 setar_hora:
tmp(381) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(382) := x"A" & "00" & '0' & x"00";	-- RET
tmp(383) := x"1" & "00" & '1' & x"41";	-- LDA R0 @SW8 AM_PM:
tmp(384) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(385) := x"7" & "00" & '1' & x"86";	-- JEQ .PM
tmp(386) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(387) := x"5" & "00" & '1' & x"01";	-- STA @LED8 R0
tmp(388) := x"5" & "00" & '0' & x"07";	-- STA @TROCA_AM_PM R0
tmp(389) := x"6" & "00" & '1' & x"89";	-- JMP .FIM_AM_PM
tmp(390) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1 PM:
tmp(391) := x"5" & "00" & '1' & x"01";	-- STA @LED8 R0
tmp(392) := x"5" & "00" & '0' & x"07";	-- STA @TROCA_AM_PM R0
tmp(393) := x"A" & "00" & '0' & x"00";	-- RET FIM_AM_PM:





		  
		  
		  
		/*
		  tmp(0) := x"9" & "00" & '0' & x"1E";	-- JSR .setup          	# Chama a função setup, para limpar os endereços
tmp(1) := x"6" & "00" & '0' & x"03";	-- JMP .LOOP_HEX
tmp(2) := x"9" & "00" & '0' & x"A6";	-- JSR .troca_hex PASSA_HEX:          # começo do LOOP para HEX0
tmp(3) := x"9" & "00" & '0' & x"4A";	-- JSR .logica_seleciona LOOP_HEX:
tmp(4) := x"7" & "00" & '0' & x"02";	-- JEQ .PASSA_HEX       	# SE botão for pressionado realiza o salto, se não continua
tmp(5) := x"9" & "00" & '0' & x"52";	-- JSR .verifica_key1
tmp(6) := x"7" & "00" & '0' & x"09";	-- JEQ .relogio_principal
tmp(7) := x"6" & "00" & '0' & x"03";	-- JMP .LOOP_HEX      	# se botão não pressionado, volta para o LOOP de HEX0
tmp(8) := x"9" & "00" & '0' & x"A3";	-- JSR .limpa_but
tmp(9) := x"9" & "00" & '0' & x"A3";	-- JSR .limpa_but relogio_principal:
tmp(10) := x"9" & "00" & '0' & x"F0";	-- JSR .verifica_carry loop_relogio:
tmp(11) := x"1" & "10" & '1' & x"41";	-- LDA R2 @SW8
tmp(12) := x"8" & "10" & '0' & x"01";	-- CEQ R2 @UM
tmp(13) := x"7" & "00" & '0' & x"13";	-- JEQ .TEMPO_RAPIDO
tmp(14) := x"4" & "11" & '0' & x"00";	-- LDI R3 $0
tmp(15) := x"5" & "11" & '1' & x"01";	-- STA @LED8 R3
tmp(16) := x"1" & "00" & '1' & x"65";	-- LDA R0 @BASE_TEMPO        		# Salva o endereço da base_tempo2 no R0
tmp(17) := x"5" & "00" & '1' & x"FD";	-- STA @LIMPA_BASE_TEMPO R0    
tmp(18) := x"6" & "00" & '0' & x"17";	-- JMP .VERIFICA_TEMPO
tmp(19) := x"4" & "11" & '0' & x"01";	-- LDI R3 $1 TEMPO_RAPIDO:
tmp(20) := x"5" & "11" & '1' & x"01";	-- STA @LED8 R3
tmp(21) := x"1" & "00" & '1' & x"66";	-- LDA R0 @BASE_TEMPO_RAP        		# Salva o endereço da base_tempo2 no R0
tmp(22) := x"5" & "00" & '1' & x"FC";	-- STA @LIMPA_BASE_TEMPO_RAP R0  
tmp(23) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM                  	# Verifica se a base de tempo será utilizada VERIFICA_TEMPO:
tmp(24) := x"7" & "00" & '0' & x"1A";	-- JEQ .INCREMENTA             	# Se for vai para a rotina de incremento
tmp(25) := x"6" & "00" & '0' & x"0A";	-- JMP .loop_relogio
tmp(26) := x"1" & "01" & '0' & x"14";	-- LDA R1 @VALOR_ATUAL0 INCREMENTA:
tmp(27) := x"2" & "01" & '0' & x"01";	-- SOMA R1 @UM
tmp(28) := x"5" & "01" & '0' & x"14";	-- STA @VALOR_ATUAL0 R1
tmp(29) := x"6" & "00" & '0' & x"0A";	-- JMP .loop_relogio
tmp(30) := x"0" & "00" & '0' & x"00";	-- NOP setup:              # Definindo a função setup, roda sempre no início limpando os valores
tmp(31) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0           
tmp(32) := x"5" & "00" & '0' & x"00";	-- STA @ZERO R0
tmp(33) := x"5" & "00" & '0' & x"06";	-- STA @ATUAL R0
tmp(34) := x"5" & "00" & '1' & x"20";	-- STA @HEX0 R0
tmp(35) := x"5" & "00" & '1' & x"21";	-- STA @HEX1 R0
tmp(36) := x"5" & "00" & '1' & x"22";	-- STA @HEX2 R0
tmp(37) := x"5" & "00" & '1' & x"23";	-- STA @HEX3 R0
tmp(38) := x"5" & "00" & '1' & x"24";	-- STA @HEX4 R0
tmp(39) := x"5" & "00" & '1' & x"25";	-- STA @HEX5 R0
tmp(40) := x"5" & "00" & '1' & x"01";	-- STA @LED8 R0
tmp(41) := x"5" & "00" & '1' & x"02";	-- STA @LED9 R0
tmp(42) := x"5" & "00" & '0' & x"0A";	-- STA @DESPERTADOR_HEX0 R0
tmp(43) := x"5" & "00" & '0' & x"0B";	-- STA @DESPERTADOR_HEX1 R0
tmp(44) := x"5" & "00" & '0' & x"0C";	-- STA @DESPERTADOR_HEX2 R0
tmp(45) := x"5" & "00" & '0' & x"0D";	-- STA @DESPERTADOR_HEX3 R0
tmp(46) := x"5" & "00" & '0' & x"0E";	-- STA @DESPERTADOR_HEX4 R0
tmp(47) := x"5" & "00" & '0' & x"0F";	-- STA @DESPERTADOR_HEX5 R0
tmp(48) := x"5" & "00" & '0' & x"14";	-- STA @VALOR_ATUAL0 R0
tmp(49) := x"5" & "00" & '0' & x"15";	-- STA @VALOR_ATUAL1 R0
tmp(50) := x"5" & "00" & '0' & x"16";	-- STA @VALOR_ATUAL2 R0
tmp(51) := x"5" & "00" & '0' & x"17";	-- STA @VALOR_ATUAL3 R0
tmp(52) := x"5" & "00" & '0' & x"18";	-- STA @VALOR_ATUAL4 R0
tmp(53) := x"5" & "00" & '0' & x"19";	-- STA @VALOR_ATUAL5 R0
tmp(54) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1
tmp(55) := x"5" & "00" & '0' & x"01";	-- STA @UM R0
tmp(56) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(57) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(58) := x"5" & "00" & '1' & x"FF";	-- STA @LIMPA_KEY0 R0
tmp(59) := x"4" & "00" & '0' & x"02";	-- LDI R0 $2
tmp(60) := x"5" & "00" & '0' & x"02";	-- STA @DOIS R0
tmp(61) := x"4" & "00" & '0' & x"03";	-- LDI R0 $3
tmp(62) := x"5" & "00" & '0' & x"03";	-- STA @TRES R0
tmp(63) := x"4" & "00" & '0' & x"04";	-- LDI R0 $4
tmp(64) := x"5" & "00" & '0' & x"04";	-- STA @QUATRO R0
tmp(65) := x"4" & "00" & '0' & x"05";	-- LDI R0 $5
tmp(66) := x"5" & "00" & '0' & x"05";	-- STA @CINCO R0
tmp(67) := x"4" & "00" & '0' & x"06";	-- LDI R0 $6
tmp(68) := x"5" & "00" & '0' & x"25";	-- STA @SEIS R0
tmp(69) := x"4" & "00" & '0' & x"0A";	-- LDI R0 $10
tmp(70) := x"5" & "00" & '0' & x"26";	-- STA @DEZ R0
tmp(71) := x"4" & "00" & '0' & x"20";	-- LDI R0 $32
tmp(72) := x"5" & "00" & '0' & x"09";	-- STA @LIMITE_LED R0
tmp(73) := x"A" & "00" & '0' & x"00";	-- RET
tmp(74) := x"9" & "00" & '0' & x"56";	-- JSR .escreveSW      	# Função que realiza a leitura e faz verificação em qual HEX está escrevendo e escreve no correto logica_seleciona:
tmp(75) := x"9" & "00" & '0' & x"E5";	-- JSR .verifica_SW9   	# Função que faz a verificação se o SW9 está ativo, se sim será 12H
tmp(76) := x"9" & "00" & '0' & x"4E";	-- JSR .verifica_key0  	# Função que faz a verificação se o botão KEY0 foi pressionado, se sim flag EQUAL = 1
tmp(77) := x"A" & "00" & '0' & x"00";	-- RET
tmp(78) := x"0" & "00" & '0' & x"00";	-- NOP verifica_key0:      # Definindo a função para verificar KEY0
tmp(79) := x"1" & "10" & '1' & x"60";	-- LDA R2 @KEY0
tmp(80) := x"8" & "10" & '0' & x"01";	-- CEQ R2 @UM
tmp(81) := x"A" & "00" & '0' & x"00";	-- RET
tmp(82) := x"0" & "00" & '0' & x"00";	-- NOP verifica_key1:      # Definindo a função para verificar KEY0
tmp(83) := x"1" & "11" & '1' & x"61";	-- LDA R3 @KEY1
tmp(84) := x"8" & "11" & '0' & x"01";	-- CEQ R3 @UM
tmp(85) := x"A" & "00" & '0' & x"00";	-- RET
tmp(86) := x"9" & "00" & '0' & x"B8";	-- JSR .VALIDA_ENTRADA escreveSW:
tmp(87) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7
tmp(88) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(89) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(90) := x"7" & "00" & '0' & x"6A";	-- JEQ .HEX0 
tmp(91) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(92) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(93) := x"7" & "00" & '0' & x"70";	-- JEQ .HEX1
tmp(94) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(95) := x"8" & "00" & '0' & x"02";	-- CEQ R0 @DOIS
tmp(96) := x"7" & "00" & '0' & x"76";	-- JEQ .HEX2 
tmp(97) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(98) := x"8" & "00" & '0' & x"03";	-- CEQ R0 @TRES
tmp(99) := x"7" & "00" & '0' & x"7C";	-- JEQ .HEX3
tmp(100) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(101) := x"8" & "00" & '0' & x"04";	-- CEQ R0 @QUATRO
tmp(102) := x"7" & "00" & '0' & x"82";	-- JEQ .HEX4
tmp(103) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(104) := x"8" & "00" & '0' & x"05";	-- CEQ R0 @CINCO
tmp(105) := x"7" & "00" & '0' & x"8E";	-- JEQ .HEX5
tmp(106) := x"1" & "00" & '0' & x"20";	-- LDA R0 @FLAG_9 HEX0:
tmp(107) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(108) := x"7" & "00" & '0' & x"99";	-- JEQ .FINAL
tmp(109) := x"5" & "01" & '1' & x"20";	-- STA @HEX0 R1
tmp(110) := x"5" & "01" & '0' & x"14";	-- STA @VALOR_ATUAL0 R1 
tmp(111) := x"6" & "00" & '0' & x"99";	-- JMP .FINAL 
tmp(112) := x"1" & "00" & '0' & x"21";	-- LDA R0 @FLAG_5 HEX1:
tmp(113) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(114) := x"7" & "00" & '0' & x"99";	-- JEQ .FINAL
tmp(115) := x"5" & "01" & '1' & x"21";	-- STA @HEX1 R1 
tmp(116) := x"5" & "01" & '0' & x"15";	-- STA @VALOR_ATUAL1 R1 
tmp(117) := x"6" & "00" & '0' & x"99";	-- JMP .FINAL 
tmp(118) := x"1" & "00" & '0' & x"20";	-- LDA R0 @FLAG_9 HEX2:
tmp(119) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(120) := x"7" & "00" & '0' & x"99";	-- JEQ .FINAL
tmp(121) := x"5" & "01" & '1' & x"22";	-- STA @HEX2 R1 
tmp(122) := x"5" & "01" & '0' & x"16";	-- STA @VALOR_ATUAL2 R1 
tmp(123) := x"6" & "00" & '0' & x"99";	-- JMP .FINAL 
tmp(124) := x"1" & "00" & '0' & x"21";	-- LDA R0 @FLAG_5 HEX3:
tmp(125) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(126) := x"7" & "00" & '0' & x"99";	-- JEQ .FINAL
tmp(127) := x"5" & "01" & '1' & x"23";	-- STA @HEX3 R1 
tmp(128) := x"5" & "01" & '0' & x"17";	-- STA @VALOR_ATUAL3 R1 
tmp(129) := x"6" & "00" & '0' & x"99";	-- JMP .FINAL 
tmp(130) := x"1" & "00" & '0' & x"1F";	-- LDA R0 @FLAG_12_OU_24 HEX4:
tmp(131) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(132) := x"7" & "00" & '0' & x"88";	-- JEQ .12_VERIFICA
tmp(133) := x"1" & "00" & '0' & x"24";	-- LDA R0 @FLAG_4
tmp(134) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(135) := x"7" & "00" & '0' & x"8B";	-- JEQ .CARREGA_HEX4
tmp(136) := x"1" & "00" & '0' & x"23";	-- LDA R0 @FLAG_2 12_VERIFICA:
tmp(137) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(138) := x"7" & "00" & '0' & x"99";	-- JEQ .FINAL
tmp(139) := x"5" & "01" & '1' & x"24";	-- STA @HEX4 R1  CARREGA_HEX4:
tmp(140) := x"5" & "01" & '0' & x"18";	-- STA @VALOR_ATUAL4 R1 
tmp(141) := x"6" & "00" & '0' & x"99";	-- JMP .FINAL 
tmp(142) := x"1" & "00" & '0' & x"1F";	-- LDA R0 @FLAG_12_OU_24 HEX5:
tmp(143) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(144) := x"7" & "00" & '0' & x"94";	-- JEQ .12_VERIFICA_5
tmp(145) := x"1" & "00" & '0' & x"23";	-- LDA R0 @FLAG_2
tmp(146) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(147) := x"7" & "00" & '0' & x"97";	-- JEQ .CARREGA_HEX5
tmp(148) := x"1" & "00" & '0' & x"22";	-- LDA R0 @FLAG_1 12_VERIFICA_5:
tmp(149) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(150) := x"7" & "00" & '0' & x"99";	-- JEQ .FINAL
tmp(151) := x"5" & "01" & '1' & x"25";	-- STA @HEX5 R1  CARREGA_HEX5:
tmp(152) := x"5" & "01" & '0' & x"19";	-- STA @VALOR_ATUAL5 R1 
tmp(153) := x"A" & "00" & '0' & x"00";	-- RET  FINAL:
tmp(154) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL atualiza_atual:
tmp(155) := x"8" & "00" & '0' & x"05";	-- CEQ R0 @CINCO
tmp(156) := x"7" & "00" & '0' & x"A0";	-- JEQ .VOLTA_UM
tmp(157) := x"2" & "00" & '0' & x"01";	-- SOMA R0 @UM
tmp(158) := x"5" & "00" & '0' & x"06";	-- STA @ATUAL R0
tmp(159) := x"A" & "00" & '0' & x"00";	-- RET
tmp(160) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0 VOLTA_UM:
tmp(161) := x"5" & "00" & '0' & x"06";	-- STA @ATUAL R0
tmp(162) := x"A" & "00" & '0' & x"00";	-- RET
tmp(163) := x"5" & "00" & '1' & x"FF";	-- STA @LIMPA_KEY0 R0  limpa_but:
tmp(164) := x"5" & "00" & '1' & x"FE";	-- STA @LIMPA_KEY1 R0
tmp(165) := x"A" & "00" & '0' & x"00";	-- RET
tmp(166) := x"9" & "00" & '0' & x"9A";	-- JSR .atualiza_atual troca_hex:
tmp(167) := x"9" & "00" & '0' & x"AB";	-- JSR .ajusta_leds
tmp(168) := x"9" & "00" & '0' & x"B5";	-- JSR .muda_led
tmp(169) := x"9" & "00" & '0' & x"A3";	-- JSR .limpa_but
tmp(170) := x"A" & "00" & '0' & x"00";	-- RET
tmp(171) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED ajusta_leds:
tmp(172) := x"8" & "00" & '0' & x"09";	-- CEQ R0 @LIMITE_LED
tmp(173) := x"7" & "00" & '0' & x"B2";	-- JEQ .VOLTA_LED
tmp(174) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(175) := x"2" & "00" & '0' & x"08";	-- SOMA R0 @AUX_LED
tmp(176) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(177) := x"A" & "00" & '0' & x"00";	-- RET
tmp(178) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1 VOLTA_LED:
tmp(179) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(180) := x"A" & "00" & '0' & x"00";	-- RET
tmp(181) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED muda_led:
tmp(182) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(183) := x"A" & "00" & '0' & x"00";	-- RET
tmp(184) := x"4" & "11" & '0' & x"01";	-- LDI R3 $1 VALIDA_ENTRADA:
tmp(185) := x"1" & "01" & '0' & x"1F";	-- LDA R1 @FLAG_12_OU_24
tmp(186) := x"8" & "01" & '0' & x"01";	-- CEQ R1 @UM 
tmp(187) := x"7" & "00" & '0' & x"C9";	-- JEQ .12H            	# Salta se estiver no modo 12HORAS se não continua para 24horas
tmp(188) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7
tmp(189) := x"C" & "01" & '0' & x"03";	-- CLT R1 @TRES
tmp(190) := x"D" & "00" & '0' & x"DF";	-- JLT .MENOR_TRES     	# modo 24 horas, verifica se o valor é menor que 3 (para validar a hora mais significativa)
tmp(191) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0           
tmp(192) := x"5" & "00" & '0' & x"23";	-- STA @FLAG_2 R0      	# desativa a escrita se a hora não é permitida
tmp(193) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7
tmp(194) := x"C" & "01" & '0' & x"05";	-- CLT R1 @CINCO
tmp(195) := x"D" & "00" & '0' & x"C7";	-- JLT .MENOR_QUATRO   	# modo 24 horas, verifica se o valor é menor que 3 (para validar a segunda hora mais significativa)
tmp(196) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(197) := x"5" & "00" & '0' & x"24";	-- STA @FLAG_4 R0      	# desativa a escrita se a hora não é permitida
tmp(198) := x"6" & "00" & '0' & x"D3";	-- JMP .COMUM
tmp(199) := x"5" & "11" & '0' & x"24";	-- STA @FLAG_4 R3  MENOR_QUATRO:
tmp(200) := x"6" & "00" & '0' & x"E0";	-- JMP .MENOR_SEIS
tmp(201) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7 12H:            # Faz a verificação no caso de 12H
tmp(202) := x"C" & "01" & '0' & x"02";	-- CLT R1 @DOIS
tmp(203) := x"D" & "00" & '0' & x"DE";	-- JLT .MENOR_DOIS         	# verifica se é menor que 2
tmp(204) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(205) := x"5" & "00" & '0' & x"22";	-- STA @FLAG_1 R0
tmp(206) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7
tmp(207) := x"C" & "01" & '0' & x"03";	-- CLT R1 @TRES
tmp(208) := x"D" & "00" & '0' & x"DF";	-- JLT .MENOR_TRES         	# verifica se é menor que 3
tmp(209) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(210) := x"5" & "00" & '0' & x"23";	-- STA @FLAG_2 R0
tmp(211) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7 COMUM:
tmp(212) := x"C" & "01" & '0' & x"25";	-- CLT R1 @SEIS
tmp(213) := x"D" & "00" & '0' & x"E0";	-- JLT .MENOR_SEIS         	# verifica se é menor que 6
tmp(214) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(215) := x"5" & "00" & '0' & x"21";	-- STA @FLAG_5 R0
tmp(216) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7
tmp(217) := x"C" & "01" & '0' & x"26";	-- CLT R1 @DEZ
tmp(218) := x"D" & "00" & '0' & x"E1";	-- JLT .MENOR_DEZ         	# verifica se é menor que 6
tmp(219) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(220) := x"5" & "00" & '0' & x"20";	-- STA @FLAG_9 R0
tmp(221) := x"6" & "00" & '0' & x"E4";	-- JMP .FINAL_FUNC
tmp(222) := x"5" & "11" & '0' & x"22";	-- STA @FLAG_1 R3      	# ATIVA SÓ QUANDO MENOR QUE 2 MENOR_DOIS: 
tmp(223) := x"5" & "11" & '0' & x"23";	-- STA @FLAG_2 R3      	# ATIVA QUANDO FOR MENOR QUE 3 MENOR_TRES:
tmp(224) := x"5" & "11" & '0' & x"21";	-- STA @FLAG_5 R3   MENOR_SEIS:
tmp(225) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1 MENOR_DEZ:
tmp(226) := x"5" & "11" & '0' & x"20";	-- STA @FLAG_9 R3  
tmp(227) := x"6" & "00" & '0' & x"E4";	-- JMP .FINAL_FUNC
tmp(228) := x"A" & "00" & '0' & x"00";	-- RET FINAL_FUNC:
tmp(229) := x"1" & "00" & '1' & x"42";	-- LDA R0 @SW9 verifica_SW9:
tmp(230) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(231) := x"7" & "00" & '0' & x"EC";	-- JEQ .SW_ATIVO
tmp(232) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0
tmp(233) := x"5" & "00" & '0' & x"1F";	-- STA @FLAG_12_OU_24 R0 
tmp(234) := x"5" & "00" & '1' & x"02";	-- STA @LED9 R0
tmp(235) := x"A" & "00" & '0' & x"00";	-- RET
tmp(236) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1 SW_ATIVO:
tmp(237) := x"5" & "00" & '0' & x"1F";	-- STA @FLAG_12_OU_24 R0 
tmp(238) := x"5" & "00" & '1' & x"02";	-- STA @LED9 R0
tmp(239) := x"A" & "00" & '0' & x"00";	-- RET
tmp(240) := x"1" & "01" & '0' & x"01";	-- LDA R1 @UM                   		# Carrega 1 no registrador para acender o LED9 verifica_carry:
tmp(241) := x"5" & "01" & '1' & x"02";	-- STA @LED9 R1                		# Acende o LED
tmp(242) := x"1" & "10" & '0' & x"14";	-- LDA R2 @VALOR_ATUAL0            	# LEITURA DE HEX0 
tmp(243) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ                     	# VERIFICA SE É IGUAL A 10 PARA O CARRY
tmp(244) := x"7" & "00" & '0' & x"F8";	-- JEQ .CARRY_DEZ_SEG              	# SALTA SE TIVER O CARRY
tmp(245) := x"1" & "10" & '0' & x"14";	-- LDA R2 @VALOR_ATUAL0            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX0
tmp(246) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(247) := x"A" & "00" & '0' & x"00";	-- RET
tmp(248) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO                    	# COMO TEVE O CARRY, ESCREVE 0 EM SEGUNDO CARRY_DEZ_SEG:
tmp(249) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(250) := x"5" & "10" & '0' & x"14";	-- STA @VALOR_ATUAL0 R2        	# ESCREVE 0 NOS SEGUNDOS QUANDO CARRY
tmp(251) := x"1" & "10" & '0' & x"15";	-- LDA R2 @VALOR_ATUAL1        	# LEITURA DO HEX1
tmp(252) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(253) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2
tmp(254) := x"8" & "10" & '0' & x"25";	-- CEQ R2 @SEIS                	# VERIFICA SE NÃO VAI TER O CARRY
tmp(255) := x"7" & "00" & '1' & x"03";	-- JEQ .CARRY_MIN              	# SALTA SE TIVER CARRY
tmp(256) := x"1" & "10" & '0' & x"15";	-- LDA R2 @VALOR_ATUAL1            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX1
tmp(257) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(258) := x"A" & "00" & '0' & x"00";	-- RET
tmp(259) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO                	# COMO TEVE CARRY ESCREVE 0 EM HEX1 CARRY_MIN:
tmp(260) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(261) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2 
tmp(262) := x"1" & "10" & '0' & x"16";	-- LDA R2 @VALOR_ATUAL2        	# LEITURA DO HEX2 PARA VER SE VAI TER CARRY
tmp(263) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(264) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2
tmp(265) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ
tmp(266) := x"7" & "00" & '1' & x"0E";	-- JEQ .CARRY_DEZ_MIN          	# SE TIVER CARRY REALIZA O SALTO
tmp(267) := x"1" & "10" & '0' & x"16";	-- LDA R2 @VALOR_ATUAL2            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX2
tmp(268) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(269) := x"A" & "00" & '0' & x"00";	-- RET
tmp(270) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO               	# COMO TEVE CARRY ESCREVE 0 EM HEX2 CARRY_DEZ_MIN:
tmp(271) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(272) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2 
tmp(273) := x"1" & "10" & '0' & x"17";	-- LDA R2 @VALOR_ATUAL3
tmp(274) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(275) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2
tmp(276) := x"8" & "10" & '0' & x"25";	-- CEQ R2 @SEIS
tmp(277) := x"7" & "00" & '1' & x"19";	-- JEQ .CARRY_HORA
tmp(278) := x"1" & "10" & '0' & x"17";	-- LDA R2 @VALOR_ATUAL3            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX3
tmp(279) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(280) := x"A" & "00" & '0' & x"00";	-- RET
tmp(281) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO CARRY_HORA:
tmp(282) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(283) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2 
tmp(284) := x"1" & "11" & '0' & x"1F";	-- LDA R3 @FLAG_12_OU_24
tmp(285) := x"8" & "11" & '0' & x"01";	-- CEQ R3 @UM
tmp(286) := x"7" & "00" & '1' & x"4D";	-- JEQ .HORA_12        	#SALTA SE O MODO DE 12 HORAS ESTIVER ATIVADO 
tmp(287) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4        	# COMEÇA A VERIFICAÇÃO PARA 24HORAS
tmp(288) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(289) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(290) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5        	# PEGA O VALOR DA HORA PARA SABER QUAL COMPARAÇÃO VOCÊ VAI FAZER
tmp(291) := x"8" & "10" & '0' & x"02";	-- CEQ R2 @DOIS 
tmp(292) := x"7" & "00" & '1' & x"2B";	-- JEQ .DEPOIS_DAS_20H
tmp(293) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(294) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ
tmp(295) := x"7" & "00" & '1' & x"45";	-- JEQ .CARRY_HORA_24
tmp(296) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX2
tmp(297) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(298) := x"A" & "00" & '0' & x"00";	-- RET                           	# ROTINA ANTES DAS 20H
tmp(299) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4 DEPOIS_DAS_20H:
tmp(300) := x"8" & "10" & '0' & x"04";	-- CEQ R2 @QUATRO 
tmp(301) := x"7" & "00" & '1' & x"37";	-- JEQ .RESET_24_HORA
tmp(302) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(303) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2 
tmp(304) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(305) := x"A" & "00" & '0' & x"00";	-- RET
tmp(306) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	#QUANDO ESTAMOS EM 20HORAS MAIS
tmp(307) := x"8" & "10" & '0' & x"04";	-- CEQ R2 @QUATRO
tmp(308) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX4 JEQ .RESET_24_HORA:
tmp(309) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(310) := x"A" & "00" & '0' & x"00";	-- RET
tmp(311) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO RESET_24_HORA:
tmp(312) := x"5" & "10" & '0' & x"14";	-- STA @VALOR_ATUAL0 R2 
tmp(313) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(314) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2 
tmp(315) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(316) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2 
tmp(317) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(318) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2
tmp(319) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(320) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(321) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(322) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(323) := x"5" & "10" & '1' & x"25";	-- STA @HEX5 R2
tmp(324) := x"A" & "00" & '0' & x"00";	-- RET
tmp(325) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO CARRY_HORA_24:
tmp(326) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(327) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2 
tmp(328) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5
tmp(329) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(330) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(331) := x"5" & "10" & '1' & x"25";	-- STA @ HEX5 R2
tmp(332) := x"A" & "00" & '0' & x"00";	-- RET
tmp(333) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4        	# LEITURA DE HEX4 HORA_12:
tmp(334) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(335) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(336) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5
tmp(337) := x"8" & "10" & '0' & x"01";	-- CEQ R2 @UM
tmp(338) := x"7" & "00" & '1' & x"59";	-- JEQ .10H_MAIS
tmp(339) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(340) := x"8" & "10" & '0' & x"26";	-- CEQ R2 @DEZ
tmp(341) := x"7" & "00" & '1' & x"63";	-- JEQ .CARRY_DEZ_HORA_12
tmp(342) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(343) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(344) := x"A" & "00" & '0' & x"00";	-- RET 
tmp(345) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4 10H_MAIS:
tmp(346) := x"8" & "10" & '0' & x"03";	-- CEQ R2 @TRES
tmp(347) := x"7" & "00" & '1' & x"6B";	-- JEQ .RESET_12H_TROCA_AM_PM
tmp(348) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4
tmp(349) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(350) := x"A" & "00" & '0' & x"00";	-- RET 
tmp(351) := x"7" & "00" & '1' & x"63";	-- JEQ .CARRY_DEZ_HORA_12
tmp(352) := x"1" & "10" & '0' & x"18";	-- LDA R2 @VALOR_ATUAL4            	# SE NÃO ESCREVE O VALOR ATUAL EM HEX2
tmp(353) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(354) := x"A" & "00" & '0' & x"00";	-- RET
tmp(355) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO CARRY_DEZ_HORA_12:
tmp(356) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2 
tmp(357) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(358) := x"1" & "10" & '0' & x"19";	-- LDA R2 @VALOR_ATUAL5
tmp(359) := x"2" & "10" & '0' & x"01";	-- SOMA R2 @UM
tmp(360) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(361) := x"5" & "10" & '1' & x"25";	-- STA @HEX5 R2
tmp(362) := x"A" & "00" & '0' & x"00";	-- RET
tmp(363) := x"1" & "10" & '0' & x"00";	-- LDA R2 @ZERO RESET_12H_TROCA_AM_PM:
tmp(364) := x"5" & "10" & '0' & x"14";	-- STA @VALOR_ATUAL0 R2 
tmp(365) := x"5" & "10" & '1' & x"20";	-- STA @HEX0 R2
tmp(366) := x"5" & "10" & '0' & x"15";	-- STA @VALOR_ATUAL1 R2 
tmp(367) := x"5" & "10" & '1' & x"21";	-- STA @HEX1 R2
tmp(368) := x"5" & "10" & '0' & x"16";	-- STA @VALOR_ATUAL2 R2 
tmp(369) := x"5" & "10" & '1' & x"22";	-- STA @HEX2 R2
tmp(370) := x"5" & "10" & '0' & x"17";	-- STA @VALOR_ATUAL3 R2
tmp(371) := x"5" & "10" & '1' & x"23";	-- STA @HEX3 R2
tmp(372) := x"5" & "10" & '0' & x"19";	-- STA @VALOR_ATUAL5 R2
tmp(373) := x"5" & "10" & '1' & x"25";	-- STA @HEX5 R2
tmp(374) := x"1" & "10" & '0' & x"01";	-- LDA R2 @UM 
tmp(375) := x"5" & "10" & '0' & x"18";	-- STA @VALOR_ATUAL4 R2
tmp(376) := x"5" & "10" & '1' & x"24";	-- STA @HEX4 R2
tmp(377) := x"A" & "00" & '0' & x"00";	-- RET
*/







		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  /*
		  tmp(0) := x"9" & "00" & '0' & x"06";	-- JSR .setup          	# Chama a função setup, para limpar os endereços
tmp(1) := x"6" & "00" & '0' & x"03";	-- JMP .LOOP_HEX
tmp(2) := x"9" & "00" & '0' & x"6B";	-- JSR .troca_hex PASSA_HEX:          # começo do LOOP para HEX0
tmp(3) := x"9" & "00" & '0' & x"2E";	-- JSR .logica_seleciona LOOP_HEX:
tmp(4) := x"7" & "00" & '0' & x"02";	-- JEQ .PASSA_HEX       	# SE botão for pressionado realiza o salto, se não continua
tmp(5) := x"6" & "00" & '0' & x"03";	-- JMP .LOOP_HEX      	# se botão não pressionado, volta para o LOOP de HEX0
tmp(6) := x"0" & "00" & '0' & x"00";	-- NOP setup:              # Definindo a função setup, roda sempre no início limpando os valores
tmp(7) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0           
tmp(8) := x"5" & "00" & '0' & x"00";	-- STA @ZERO R0
tmp(9) := x"5" & "00" & '0' & x"06";	-- STA @ATUAL R0
tmp(10) := x"5" & "00" & '1' & x"20";	-- STA @HEX0 R0
tmp(11) := x"5" & "00" & '1' & x"21";	-- STA @HEX1 R0
tmp(12) := x"5" & "00" & '1' & x"22";	-- STA @HEX2 R0
tmp(13) := x"5" & "00" & '1' & x"23";	-- STA @HEX3 R0
tmp(14) := x"5" & "00" & '1' & x"24";	-- STA @HEX4 R0
tmp(15) := x"5" & "00" & '1' & x"25";	-- STA @HEX5 R0
tmp(16) := x"5" & "00" & '1' & x"01";	-- STA @LED8 R0
tmp(17) := x"5" & "00" & '1' & x"02";	-- STA @LED9 R0
tmp(18) := x"5" & "00" & '0' & x"0A";	-- STA @DESPERTADOR_HEX0 R0
tmp(19) := x"5" & "00" & '0' & x"0B";	-- STA @DESPERTADOR_HEX1 R0
tmp(20) := x"5" & "00" & '0' & x"0C";	-- STA @DESPERTADOR_HEX2 R0
tmp(21) := x"5" & "00" & '0' & x"0D";	-- STA @DESPERTADOR_HEX3 R0
tmp(22) := x"5" & "00" & '0' & x"0E";	-- STA @DESPERTADOR_HEX4 R0
tmp(23) := x"5" & "00" & '0' & x"0F";	-- STA @DESPERTADOR_HEX5 R0
tmp(24) := x"5" & "00" & '0' & x"14";	-- STA @VALOR_ATUAL0 R0
tmp(25) := x"5" & "00" & '0' & x"15";	-- STA @VALOR_ATUAL1 R0
tmp(26) := x"5" & "00" & '0' & x"16";	-- STA @VALOR_ATUAL2 R0
tmp(27) := x"5" & "00" & '0' & x"17";	-- STA @VALOR_ATUAL3 R0
tmp(28) := x"5" & "00" & '0' & x"18";	-- STA @VALOR_ATUAL4 R0
tmp(29) := x"5" & "00" & '0' & x"19";	-- STA @VALOR_ATUAL5 R0
tmp(30) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1
tmp(31) := x"5" & "00" & '0' & x"01";	-- STA @UM R0
tmp(32) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(33) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(34) := x"5" & "00" & '1' & x"FF";	-- STA @LIMPA_KEY0 R0
tmp(35) := x"4" & "00" & '0' & x"02";	-- LDI R0 $2
tmp(36) := x"5" & "00" & '0' & x"02";	-- STA @DOIS R0
tmp(37) := x"4" & "00" & '0' & x"03";	-- LDI R0 $3
tmp(38) := x"5" & "00" & '0' & x"03";	-- STA @TRES R0
tmp(39) := x"4" & "00" & '0' & x"04";	-- LDI R0 $4
tmp(40) := x"5" & "00" & '0' & x"04";	-- STA @QUATRO R0
tmp(41) := x"4" & "00" & '0' & x"05";	-- LDI R0 $5
tmp(42) := x"5" & "00" & '0' & x"05";	-- STA @CINCO R0
tmp(43) := x"4" & "00" & '0' & x"20";	-- LDI R0 $32
tmp(44) := x"5" & "00" & '0' & x"09";	-- STA @LIMITE_LED R0
tmp(45) := x"A" & "00" & '0' & x"00";	-- RET
tmp(46) := x"9" & "00" & '0' & x"35";	-- JSR .escreveSW      	# Função que realiza a leitura e faz verificação em qual HEX está escrevendo e escreve no correto logica_seleciona:
tmp(47) := x"9" & "00" & '0' & x"31";	-- JSR .verifica_key0  	# Função que faz a verificação se o botão KEY0 foi pressionado, se sim flag EQUAL = 1
tmp(48) := x"A" & "00" & '0' & x"00";	-- RET
tmp(49) := x"0" & "00" & '0' & x"00";	-- NOP verifica_key0:      # Definindo a função para verificar KEY0
tmp(50) := x"1" & "10" & '1' & x"60";	-- LDA R2 @KEY0
tmp(51) := x"8" & "10" & '0' & x"01";	-- CEQ R2 @UM
tmp(52) := x"A" & "00" & '0' & x"00";	-- RET
tmp(53) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7 escreveSW:
tmp(54) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(55) := x"8" & "00" & '0' & x"00";	-- CEQ R0 @ZERO
tmp(56) := x"7" & "00" & '0' & x"48";	-- JEQ .HEX0 
tmp(57) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(58) := x"8" & "00" & '0' & x"01";	-- CEQ R0 @UM
tmp(59) := x"7" & "00" & '0' & x"4B";	-- JEQ .HEX1
tmp(60) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(61) := x"8" & "00" & '0' & x"02";	-- CEQ R0 @DOIS
tmp(62) := x"7" & "00" & '0' & x"4E";	-- JEQ .HEX2 
tmp(63) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(64) := x"8" & "00" & '0' & x"03";	-- CEQ R0 @TRES
tmp(65) := x"7" & "00" & '0' & x"51";	-- JEQ .HEX3
tmp(66) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(67) := x"8" & "00" & '0' & x"04";	-- CEQ R0 @QUATRO
tmp(68) := x"7" & "00" & '0' & x"54";	-- JEQ .HEX4
tmp(69) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL
tmp(70) := x"8" & "00" & '0' & x"05";	-- CEQ R0 @CINCO
tmp(71) := x"7" & "00" & '0' & x"57";	-- JEQ .HEX5
tmp(72) := x"5" & "01" & '1' & x"20";	-- STA @HEX0 R1 HEX0:
tmp(73) := x"5" & "01" & '0' & x"14";	-- STA @VALOR_ATUAL0 R1 
tmp(74) := x"6" & "00" & '0' & x"59";	-- JMP .FINAL 
tmp(75) := x"5" & "01" & '1' & x"21";	-- STA @HEX1 R1  HEX1:
tmp(76) := x"5" & "01" & '0' & x"15";	-- STA @VALOR_ATUAL1 R1 
tmp(77) := x"6" & "00" & '0' & x"59";	-- JMP .FINAL 
tmp(78) := x"5" & "01" & '1' & x"22";	-- STA @HEX2 R1  HEX2:
tmp(79) := x"5" & "01" & '0' & x"16";	-- STA @VALOR_ATUAL2 R1 
tmp(80) := x"6" & "00" & '0' & x"59";	-- JMP .FINAL 
tmp(81) := x"5" & "01" & '1' & x"23";	-- STA @HEX3 R1  HEX3:
tmp(82) := x"5" & "01" & '0' & x"17";	-- STA @VALOR_ATUAL3 R1 
tmp(83) := x"6" & "00" & '0' & x"59";	-- JMP .FINAL 
tmp(84) := x"5" & "01" & '1' & x"24";	-- STA @HEX4 R1  HEX4:
tmp(85) := x"5" & "01" & '0' & x"18";	-- STA @VALOR_ATUAL4 R1 
tmp(86) := x"6" & "00" & '0' & x"59";	-- JMP .FINAL 
tmp(87) := x"5" & "01" & '1' & x"25";	-- STA @HEX5 R1  HEX5:
tmp(88) := x"5" & "01" & '0' & x"19";	-- STA @VALOR_ATUAL5 R1 
tmp(89) := x"A" & "00" & '0' & x"00";	-- RET  FINAL:
tmp(90) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL atualiza_atual:
tmp(91) := x"8" & "00" & '0' & x"05";	-- CEQ R0 @CINCO
tmp(92) := x"7" & "00" & '0' & x"60";	-- JEQ .VOLTA_UM
tmp(93) := x"2" & "00" & '0' & x"01";	-- SOMA R0 @UM
tmp(94) := x"5" & "00" & '0' & x"06";	-- STA @ATUAL R0
tmp(95) := x"A" & "00" & '0' & x"00";	-- RET
tmp(96) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0 VOLTA_UM:
tmp(97) := x"5" & "00" & '0' & x"06";	-- STA @ATUAL R0
tmp(98) := x"A" & "00" & '0' & x"00";	-- RET
tmp(99) := x"1" & "00" & '0' & x"06";	-- LDA R0 @ATUAL COMP_ATUAL:
tmp(100) := x"8" & "00" & '0' & x"07";	-- CEQ R0 @CONT
tmp(101) := x"9" & "00" & '0' & x"73";	-- JSR .atualiza_cont
tmp(102) := x"1" & "01" & '1' & x"40";	-- LDA R1 @SW0a7
tmp(103) := x"A" & "00" & '0' & x"00";	-- RET
tmp(104) := x"5" & "00" & '1' & x"FF";	-- STA @LIMPA_KEY0 R0  limpa_but:
tmp(105) := x"5" & "00" & '1' & x"FE";	-- STA @LIMPA_KEY1 R0
tmp(106) := x"A" & "00" & '0' & x"00";	-- RET
tmp(107) := x"9" & "00" & '0' & x"5A";	-- JSR .atualiza_atual troca_hex:
tmp(108) := x"9" & "00" & '0' & x"77";	-- JSR .ajusta_leds
tmp(109) := x"9" & "00" & '0' & x"81";	-- JSR .muda_led
tmp(110) := x"9" & "00" & '0' & x"68";	-- JSR .limpa_but
tmp(111) := x"A" & "00" & '0' & x"00";	-- RET
tmp(112) := x"4" & "00" & '0' & x"00";	-- LDI R0 $0 def_cont:
tmp(113) := x"5" & "00" & '0' & x"07";	-- STA @CONT R0
tmp(114) := x"A" & "00" & '0' & x"00";	-- RET
tmp(115) := x"1" & "00" & '0' & x"01";	-- LDA R0 @UM atualiza_cont:
tmp(116) := x"2" & "00" & '0' & x"01";	-- SOMA R0 @UM
tmp(117) := x"5" & "00" & '0' & x"07";	-- STA @CONT R0
tmp(118) := x"A" & "00" & '0' & x"00";	-- RET
tmp(119) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED ajusta_leds:
tmp(120) := x"8" & "00" & '0' & x"09";	-- CEQ R0 @LIMITE_LED
tmp(121) := x"7" & "00" & '0' & x"7E";	-- JEQ .VOLTA_LED
tmp(122) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED
tmp(123) := x"2" & "00" & '0' & x"08";	-- SOMA R0 @AUX_LED
tmp(124) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(125) := x"A" & "00" & '0' & x"00";	-- RET
tmp(126) := x"4" & "00" & '0' & x"01";	-- LDI R0 $1 VOLTA_LED:
tmp(127) := x"5" & "00" & '0' & x"08";	-- STA @AUX_LED R0
tmp(128) := x"A" & "00" & '0' & x"00";	-- RET
tmp(129) := x"1" & "00" & '0' & x"08";	-- LDA R0 @AUX_LED muda_led:
tmp(130) := x"5" & "00" & '1' & x"00";	-- STA @LED0A7 R0
tmp(131) := x"A" & "00" & '0' & x"00";	-- RET
*/











        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;